CircuitMaker Text
5.6
Probes: 1
D1_A
Operating Point
0 470 191 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
100 0 30 200 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
8
5 SAVE-
218 418 106 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3798 0 0
2
5.90005e-315 0
0
11 Multimeter~
205 251 59 0 21 21
0 3 6 7 4 0 0 0 0 0
32 51 55 48 46 54 117 65 0 0
0 86
0
0 0 16448 0
6 1.000u
-21 -19 21 -11
3 MM1
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
6884 0 0
2
5.90005e-315 0
0
11 Multimeter~
205 766 166 0 21 21
0 5 8 9 2 0 0 0 0 0
32 54 50 57 46 52 109 86 0 0
0 82
0
0 0 16448 0
8 100.0Meg
-28 -19 28 -11
3 MM0
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
4807 0 0
2
5.90005e-315 0
0
7 Ground~
168 467 298 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9591 0 0
2
5.90005e-315 0
0
8 Battery~
219 174 305 0 2 5
0 3 2
0
0 0 864 0
2 1V
16 -2 30 6
2 V1
16 -12 30 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6279 0 0
2
5.90005e-315 0
0
7 Ground~
168 174 347 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4515 0 0
2
5.90005e-315 0
0
6 Diode~
219 467 228 0 2 5
0 5 2
0
0 0 832 270
5 DIODE
11 0 46 8
2 D1
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
4396 0 0
2
5.90005e-315 0
0
11 Resistor:A~
219 471 113 0 2 5
0 5 4
0
0 0 864 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6796 0 0
2
5.90005e-315 0
0
7
1 1 3 0 0 4224 0 2 5 0 0 4
226 82
226 193
174 193
174 292
2 4 4 0 0 4224 0 8 2 0 0 3
471 95
276 95
276 82
4 0 2 0 0 8320 0 3 0 0 5 3
791 189
791 264
467 264
1 0 5 0 0 4224 0 3 0 0 6 2
741 189
471 189
2 1 2 0 0 0 0 7 4 0 0 2
467 238
467 292
1 1 5 0 0 0 0 8 7 0 0 3
471 131
471 218
467 218
2 1 2 0 0 0 0 5 6 0 0 2
174 316
174 341
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
